alu_agent.sv		  file.txt    nombre.txt    salida.txt	      test.sv
alu_env.sv		  git.sh      numeros.cpp   script	      test.txt
backup.txt		  jenkins.sh  pruebas2.cpp  sim_cov_commands  upload.sh
bash_snps_xt018-AMS_2017  leer	      pruebas.cpp   test
design.sv		  nombre      prueba.txt    testbench.sv
file			  nombre.cpp  regresion     test.cpp
