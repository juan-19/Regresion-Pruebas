alu_agent.sv		  file.txt     pruebas2.cpp	 test
alu_driver.sv		  git.sh       pruebas.cpp	 testbench.sv
alu_env.sv		  jenkins.sh   prueba.txt	 test.cpp
alu_scoreboard.sv	  leer	       README.md	 test.sv
backup.txt		  nombre       regresion	 test.txt
bash_snps_xt018-AMS_2017  nombre.cpp   salida.txt	 upload.sh
design.sv		  nombre.txt   script
file			  numeros.cpp  sim_cov_commands
