alu_env.sv		  file.txt    numeros.cpp   script	      test.txt
backup.txt		  git.sh      pruebas2.cpp  sim_cov_commands  upload.sh
bash_snps_xt018-AMS_2017  leer	      pruebas.cpp   test
config			  nombre      prueba.txt    testbench.sv
design.sv		  nombre.cpp  regresion     test.cpp
file			  nombre.txt  salida.txt    test.sv
