alu_agent.sv		  design.sv   nombre	    README.md	      test.cpp
alu_driver.sv		  dir	      nombre.cpp    regresion	      test.sv
alu_env.sv		  file	      nombre.txt    salida.txt	      test.txt
alu_interface.sv	  file.txt    numeros.cpp   script	      upload.sh
alu_monitor.sv		  git.sh      pruebas2.cpp  sim_cov_commands
backup.txt		  jenkins.sh  pruebas.cpp   test
bash_snps_xt018-AMS_2017  leer	      prueba.txt    testbench.sv
