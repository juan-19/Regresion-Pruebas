backup.txt		  nombre	prueba.txt	  testbench.sv
bash_snps_xt018-AMS_2017  nombre.cpp	regresion	  test.cpp
file			  nombre.txt	salida.txt	  test.sv
file.txt		  numeros.cpp	script		  test.txt
git.sh			  pruebas2.cpp	sim_cov_commands  upload.sh
leer			  pruebas.cpp	test
