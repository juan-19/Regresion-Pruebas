alu_env.sv		  leer		prueba.txt	  test.cpp
backup.txt		  nombre	regresion	  test.sv
bash_snps_xt018-AMS_2017  nombre.cpp	salida.txt	  test.txt
design.sv		  nombre.txt	script		  upload.sh
file			  numeros.cpp	sim_cov_commands
file.txt		  pruebas2.cpp	test
git.sh			  pruebas.cpp	testbench.sv
