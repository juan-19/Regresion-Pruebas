file  testbench.sv
