backup.txt		  git.sh      numeros.cpp   salida.txt	      test.cpp
bash_snps_xt018-AMS_2017  leer	      pruebas2.cpp  script	      test.sv
design.sv		  nombre      pruebas.cpp   sim_cov_commands  test.txt
file			  nombre.cpp  prueba.txt    test	      upload.sh
file.txt		  nombre.txt  regresion     testbench.sv
